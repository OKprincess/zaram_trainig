// ===================================================
//	=================[ VLSISYS Lab. ]=================
//	* Author		: oksj (oksj@sookmyung.ac.kr)
//	* Filename		: click_network.v
//	* Description	: 
// ===================================================
`include		"dff.v"
`include		"click.v"

module click_network 
(
	output		o_fire_IF,o_fire_ID, o_fire_EX, o_fire_MEM, o_fire_WB,
	output		
);
	
endmodule
